// TASK: Clock Generator
task automatic tsk_clock_gen(output logic i_clk, input int CLOCK_PERIOD);
  begin
    i_clk = 1'b0;
    forever #(CLOCK_PERIOD) i_clk = !i_clk;
  end
endtask

// TASK: Reset is low active for a period of "RESET_PERIOD"
task automatic tsk_reset(output logic i_reset, input int RESET_PERIOD);
  begin
    i_reset = 1'b0; // Easter Egg
    #(RESET_PERIOD);
    i_reset = 1'b1; //
  end
endtask

// TASK: Timeout, assume after a period of "TIMEOUT",
// the design is supposed to be "PASSED"
task automatic tsk_timeout(input int TIMEOUT);
  begin
    #TIMEOUT;
    $display("\nTimeout...\n");
    $finish;
  end
endtask
