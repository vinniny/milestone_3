`timescale 1ns / 1ps
// ============================================================================
// Module: tb_hexled
// Description: Testbench to verify HEXLED (7-segment display) outputs
//              Tests counter_v3.hex program with switches and displays
// ============================================================================

module tb_hexled;

  // Clock and reset
  logic        clk;
  logic        reset;
  
  // Processor debug signals
  logic [31:0] pc_frontend;
  logic [31:0] pc_commit;
  logic        insn_vld;
  logic        halt;
  logic [3:0]  model_id;
  
  // I/O signals
  logic [31:0] io_ledr;
  logic [31:0] io_ledg;
  logic [ 6:0] io_hex0, io_hex1, io_hex2, io_hex3;
  logic [ 6:0] io_hex4, io_hex5, io_hex6, io_hex7;
  logic [31:0] io_lcd;
  logic [31:0] io_sw;
  
  // Test control
  integer      cycle_count;
  integer      test_errors;
  logic [31:0] expected_hex_low;
  logic [31:0] expected_hex_high;
  
  // Counter tracking
  logic [31:0] last_counter_value;
  logic [31:0] current_counter_value;
  integer      increment_count;
  
  // Test variables
  integer      pause_checks;
  integer      pause_errors;
  integer      addr_test_errors;
  logic [3:0]  ones, tens, new_ones, new_tens;
  integer      start_cycles;
  logic [31:0] start_value, end_value, pause_value, resume_value;
  integer      elapsed_cycles, counter_delta;
  
  // 7-segment decoder for display (active-low)
  function [6:0] digit_to_7seg(input [3:0] digit);
    case (digit)
      4'd0: digit_to_7seg = 7'h40;  // 0
      4'd1: digit_to_7seg = 7'h79;  // 1
      4'd2: digit_to_7seg = 7'h24;  // 2
      4'd3: digit_to_7seg = 7'h30;  // 3
      4'd4: digit_to_7seg = 7'h19;  // 4
      4'd5: digit_to_7seg = 7'h12;  // 5
      4'd6: digit_to_7seg = 7'h02;  // 6
      4'd7: digit_to_7seg = 7'h78;  // 7
      4'd8: digit_to_7seg = 7'h00;  // 8
      4'd9: digit_to_7seg = 7'h10;  // 9
      default: digit_to_7seg = 7'h7F;  // blank
    endcase
  endfunction
  
  // DUT instantiation
  pipelined dut (
    .i_clk(clk),
    .i_reset(reset),
    .o_pc_frontend(pc_frontend),
    .o_pc_commit(pc_commit),
    .o_insn_vld(insn_vld),
    .o_halt(halt),
    .o_model_id(model_id),
    .o_ctrl(),
    .o_mispred(),
    .o_io_ledr(io_ledr),
    .o_io_ledg(io_ledg),
    .o_io_hex0(io_hex0),
    .o_io_hex1(io_hex1),
    .o_io_hex2(io_hex2),
    .o_io_hex3(io_hex3),
    .o_io_hex4(io_hex4),
    .o_io_hex5(io_hex5),
    .o_io_hex6(io_hex6),
    .o_io_hex7(io_hex7),
    .o_io_lcd(io_lcd),
    .i_io_sw(io_sw)
  );
  
  // Clock generation (100 MHz = 10ns period)
  initial begin
    clk = 0;
    forever #5 clk = ~clk;
  end
  
  // Cycle counter
  always @(posedge clk) begin
    if (~reset)
      cycle_count <= 0;
    else
      cycle_count <= cycle_count + 1;
  end
  
  // Timeout watchdog - 2s timeout
  initial begin
    $display("⏱️  Timeout watchdog started (2s limit)...");
    #2_000_000_000; // 2s = 200,000,000 cycles @ 10ns period
    $display("\n");
    $display("⚠️  ═══════════════════════════════════════════════════════════════");
    $display("⚠️  TIMEOUT: Test exceeded 2s simulation time");
    $display("⚠️  ═══════════════════════════════════════════════════════════════");
    $display("   Cycles simulated: %0d", cycle_count);
    $display("   PC at timeout: 0x%h", pc_commit);
    $display("\n   This may indicate:");
    $display("     - Delay loops are still too long");
    $display("     - Processor stuck in infinite loop");
    $display("     - Need to use counter_v3_fast.hex\n");
    $finish;
  end
  
  // Monitor task to display HEXLED values
  task display_hexleds;
    input string label;
    logic [3:0] d0, d1, d2, d3, d4, d5;
    begin
      d0 = decode_7seg(io_hex0);
      d1 = decode_7seg(io_hex1);
      d2 = decode_7seg(io_hex2);
      d3 = decode_7seg(io_hex3);
      d4 = decode_7seg(io_hex4);
      d5 = decode_7seg(io_hex5);
      
      $display("  [%s] HEX Displays:", label);
      $display("    Raw 7-seg codes:");
      $display("      HEX7-4: %h %h %h %h", io_hex7, io_hex6, io_hex5, io_hex4);
      $display("      HEX3-0: %h %h %h %h", io_hex3, io_hex2, io_hex1, io_hex0);
      $display("    Decoded digits: %0d%0d:%0d%0d:%0d%0d (MM:SS:CC)",
               d5, d4, d3, d2, d1, d0);
      $display("    Counter value: %0d", get_counter_value());
    end
  endtask
  
  // Function to decode 7-segment to digit
  function [3:0] decode_7seg(input [6:0] segments);
    case (segments)
      7'h40: decode_7seg = 4'd0;
      7'h79: decode_7seg = 4'd1;
      7'h24: decode_7seg = 4'd2;
      7'h30: decode_7seg = 4'd3;
      7'h19: decode_7seg = 4'd4;
      7'h12: decode_7seg = 4'd5;
      7'h02: decode_7seg = 4'd6;
      7'h78: decode_7seg = 4'd7;
      7'h00: decode_7seg = 4'd8;
      7'h10: decode_7seg = 4'd9;
      7'h7F: decode_7seg = 4'd15; // blank
      default: decode_7seg = 4'd15;
    endcase
  endfunction
  
  // Get current counter value from displays (as packed BCD for comparison)
  // Returns: bits[23:0] = HEX5|HEX4|HEX3|HEX2|HEX1|HEX0 (4 bits each)
  function [31:0] get_counter_value;
    logic [3:0] d0, d1, d2, d3, d4, d5;
    d0 = decode_7seg(io_hex0);
    d1 = decode_7seg(io_hex1);
    d2 = decode_7seg(io_hex2);
    d3 = decode_7seg(io_hex3);
    d4 = decode_7seg(io_hex4);
    d5 = decode_7seg(io_hex5);
    // Return as packed BCD (4 bits per digit)
    get_counter_value = {8'h0, d5[3:0], d4[3:0], d3[3:0], d2[3:0], d1[3:0], d0[3:0]};
  endfunction
  
  // Verify all digits are valid (0-9)
  function bit all_digits_valid;
    logic [3:0] d0, d1, d2, d3, d4, d5;
    d0 = decode_7seg(io_hex0);
    d1 = decode_7seg(io_hex1);
    d2 = decode_7seg(io_hex2);
    d3 = decode_7seg(io_hex3);
    d4 = decode_7seg(io_hex4);
    d5 = decode_7seg(io_hex5);
    // Valid if digit is 0-9 or 15 (blank)
    all_digits_valid = (d0 < 10 || d0 == 15) &&
                       (d1 < 10 || d1 == 15) &&
                       (d2 < 10 || d2 == 15) &&
                       (d3 < 10 || d3 == 15) &&
                       (d4 < 10 || d4 == 15) &&
                       (d5 < 10 || d5 == 15);
  endfunction
  
  // Verify BCD encoding (digits 1 and 3 should be 0-5, others 0-9)
  // Blank displays (15) are also valid
  function bit bcd_encoding_valid;
    logic [3:0] d0, d1, d2, d3, d4, d5;
    d0 = decode_7seg(io_hex0);
    d1 = decode_7seg(io_hex1);
    d2 = decode_7seg(io_hex2);
    d3 = decode_7seg(io_hex3);
    d4 = decode_7seg(io_hex4);
    d5 = decode_7seg(io_hex5);
    // Tens digits (1, 3, 5) should be 0-5 or blank (15)
    // Ones digits (0, 2, 4) should be 0-9 or blank (15)
    bcd_encoding_valid = (d1 <= 5 || d1 == 15) && (d3 <= 5 || d3 == 15) && (d5 <= 5 || d5 == 15) &&
                         (d0 <= 9 || d0 == 15) && (d2 <= 9 || d2 == 15) && (d4 <= 9 || d4 == 15);
  endfunction
  
  // Verification task
  task verify_hexled;
    input [6:0] expected_hex0;
    input [6:0] expected_hex1;
    input [6:0] expected_hex2;
    input [6:0] expected_hex3;
    input string test_name;
    begin
      if (io_hex0 !== expected_hex0 || io_hex1 !== expected_hex1 ||
          io_hex2 !== expected_hex2 || io_hex3 !== expected_hex3) begin
        $display("  ❌ FAIL: %s", test_name);
        $display("    Expected HEX3-0: %h %h %h %h", 
                 expected_hex3, expected_hex2, expected_hex1, expected_hex0);
        $display("    Got      HEX3-0: %h %h %h %h", 
                 io_hex3, io_hex2, io_hex1, io_hex0);
        test_errors = test_errors + 1;
      end else begin
        $display("  ✅ PASS: %s", test_name);
        $display("    HEX3-0 = %h %h %h %h (digits: %0d%0d:%0d%0d)", 
                 io_hex3, io_hex2, io_hex1, io_hex0,
                 decode_7seg(io_hex3), decode_7seg(io_hex2),
                 decode_7seg(io_hex1), decode_7seg(io_hex0));
      end
    end
  endtask
  
  // Task to wait for counter increment (fixed to work with BCD)
  task wait_for_increment;
    input integer max_cycles;
    input string test_desc;
    integer i;
    logic [31:0] task_start_value, curr_value;
    begin
      task_start_value = get_counter_value();
      $display("    Waiting for increment from 0x%h (max %0d cycles)...", start_value, max_cycles);
      
      for (i = 0; i < max_cycles; i = i + 1) begin
        @(posedge clk);
        curr_value = get_counter_value();
        if (curr_value != task_start_value) begin
          $display("    ✅ Counter incremented after %0d cycles", i);
          $display("    0x%h -> 0x%h", task_start_value, curr_value);
          return;
        end
      end
      
      $display("    ⚠️  WARNING: %s - No increment after %0d cycles", test_desc, max_cycles);
      $display("    Value stayed at: 0x%h", task_start_value);
    end
  endtask
  
  // Task to verify counter increment sequence (fixed for BCD wrapping)
  task verify_increment_sequence;
    input integer num_checks;
    input integer cycles_between;
    integer i;
    logic [31:0] prev_value, curr_value;
    integer errors;
    begin
      errors = 0;
      prev_value = get_counter_value();
      $display("    Starting value: 0x%h", prev_value);
      
      for (i = 0; i < num_checks; i = i + 1) begin
        repeat(cycles_between) @(posedge clk);
        curr_value = get_counter_value();
        
        // For BCD counter, any change is acceptable (wraps at 10, 100, etc)
        if (curr_value == prev_value) begin
          $display("    ⚠️  No change: 0x%h (check %0d/%0d)", curr_value, i+1, num_checks);
          errors = errors + 1;
        end else begin
          $display("    ✓ 0x%h -> 0x%h", prev_value, curr_value);
        end
        
        prev_value = curr_value;
      end
      
      if (errors == 0) begin
        $display("  ✅ PASS: Counter incremented in all checks");
      end else begin
        $display("  ❌ FAIL: %0d checks showed no increment", errors);
        test_errors = test_errors + 1;
      end
    end
  endtask
  
  // Main test sequence
  initial begin
    $display("\n");
    $display("╔══════════════════════════════════════════════════════════════════╗");
    $display("║      HEXLED In-Depth Verification Test (counter_v3.hex)         ║");
    $display("╚══════════════════════════════════════════════════════════════════╝");
    $display("");
    
    // Initialize
    reset = 0;
    io_sw = 32'h0;
    cycle_count = 0;
    test_errors = 0;
    increment_count = 0;
    
    // Reset sequence
    $display("[INIT] Applying reset...");
    #20;
    reset = 1;
    #200;  // Give enough time after reset
    $display("[INIT] Reset released, processor running");
    $display("");
    
    // Wait for processor to initialize displays
    $display("━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━");
    $display("TEST 1: Initialization & Reset Verification");
    $display("━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━");
    
    // Start with switch on (counter enabled from the start for simple version)
    io_sw = 32'h1;
    repeat(1000) @(posedge clk);
    
    display_hexleds("Initial State (SW[0]=1)");
    
    // Verify program is running and displays are initialized
    $display("  Counter program initialized");
    
    // Check if counter is incrementing (simple check)
    last_counter_value = get_counter_value();
    repeat(1000) @(posedge clk);
    current_counter_value = get_counter_value();
    
    if (current_counter_value != last_counter_value) begin
      $display("  ✅ PASS: Counter is running");
    end else begin
      $display("  ⚠️  WARNING: Counter not incrementing in first 1000 cycles");
      $display("    Value: 0x%h", current_counter_value);
    end
    $display("");
    
    // Now verify counter continues running
    $display("━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━");
    $display("TEST 2: Display Validation");
    $display("━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━");
    
    io_sw = 32'h1;  // Ensure counter is enabled
    $display("  SW[0] = 1 (counter enabled)");
    
    // Wait a bit for displays to update
    repeat(1000) @(posedge clk);
    
    display_hexleds("After Startup");
    
    // Verify all digits are valid
    if (all_digits_valid()) begin
      $display("  ✅ PASS: All HEX displays show valid digits (0-9)");
    end else begin
      $display("  ❌ FAIL: Some displays show invalid digits");
      test_errors = test_errors + 1;
    end
    $display("");
    
    // Test 3: 7-Segment Encoding Validation  
    $display("━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━");
    $display("TEST 3: 7-Segment Encoding Validation");
    $display("━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━");
    
    $display("  Current display state:");
    $display("  Digit | Expected | HEX0 | HEX1 | HEX2 | HEX3 | HEX4 | HEX5");
    $display("  ------|----------|------|------|------|------|------|------");
    
    for (int digit = 0; digit <= 9; digit++) begin
      logic [6:0] expected_code;
      logic [3:0] digit_4bit;
      digit_4bit = digit[3:0];
      expected_code = digit_to_7seg(digit_4bit);
      $display("    %0d   |   0x%h   | %s | %s | %s | %s | %s | %s",
               digit, expected_code,
               (decode_7seg(io_hex0) == digit_4bit) ? "✓" : " ",
               (decode_7seg(io_hex1) == digit_4bit) ? "✓" : " ",
               (decode_7seg(io_hex2) == digit_4bit) ? "✓" : " ",
               (decode_7seg(io_hex3) == digit_4bit) ? "✓" : " ",
               (decode_7seg(io_hex4) == digit_4bit) ? "✓" : " ",
               (decode_7seg(io_hex5) == digit_4bit) ? "✓" : " ");
    end
    
    // Verify BCD encoding constraints
    if (bcd_encoding_valid()) begin
      $display("  ✅ PASS: BCD encoding is valid (tens digits 0-5, ones digits 0-9)");
    end else begin
      $display("  ❌ FAIL: BCD encoding invalid");
      test_errors = test_errors + 1;
    end
    $display("");
    
    // Test 4: First Increment
    $display("━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━");
    $display("TEST 4: First Counter Increment");
    $display("━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━");
    
    $display("  Counter is already enabled (SW[0]=1)");
    
    last_counter_value = get_counter_value();
    $display("  Current counter value: 0x%h", last_counter_value);
    
    // Wait for first increment (with 10-cycle delay, should happen quickly)
    wait_for_increment(200, "First increment");
    
    current_counter_value = get_counter_value();
    display_hexleds("After First Increment");
    
    // For BCD, just check that value changed (any change is valid)
    if (current_counter_value != last_counter_value) begin
      $display("  ✅ PASS: Counter incremented (0x%h -> 0x%h)", 
               last_counter_value, current_counter_value);
      increment_count = increment_count + 1;
    end else begin
      $display("  ❌ FAIL: Counter did not increment");
      test_errors = test_errors + 1;
    end
    
    // Verify digits are still valid
    if (all_digits_valid()) begin
      $display("  ✅ PASS: All digits valid after increment");
    end else begin
      $display("  ❌ FAIL: Invalid digits detected");
      test_errors = test_errors + 1;
    end
    $display("");
    
    // Test 5: Multiple Increment Sequence
    $display("━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━");
    $display("TEST 5: Multiple Increment Sequence");
    $display("━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━");
    
    $display("  Checking 5 consecutive increments (200 cycles between checks)...");
    verify_increment_sequence(5, 200);
    $display("");
    
    // Test 6: Pause Functionality
    $display("━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━");
    $display("TEST 6: Pause Functionality (SW[0] = 0)");
    $display("━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━");
    
    io_sw = 32'h0;  // Clear SW[0] to pause
    $display("  SW[0] = 0 (counter paused)");
    
    last_counter_value = get_counter_value();
    display_hexleds("At pause");
    
    // Wait a bit for any in-flight instructions to complete
    repeat(100) @(posedge clk);
    last_counter_value = get_counter_value();  // Get settled value
    
    // Wait and check multiple times to ensure it stays paused
    pause_checks = 3;
    pause_errors = 0;
    
    for (int i = 0; i < pause_checks; i++) begin
      repeat(1000) @(posedge clk);  // Wait longer to ensure no change
      current_counter_value = get_counter_value();
      
      if (current_counter_value != last_counter_value) begin
        $display("  ❌ Check %0d: Counter changed while paused (0x%h -> 0x%h)", 
                 i+1, last_counter_value, current_counter_value);
        pause_errors = pause_errors + 1;
        last_counter_value = current_counter_value;  // Update for next check
      end else begin
        $display("  ✓ Check %0d: Counter stable at 0x%h", i+1, current_counter_value);
      end
    end
    
    if (pause_errors == 0) begin
      $display("  ✅ PASS: Counter correctly paused (verified %0d times)", pause_checks);
    end else begin
      $display("  ⚠️  WARNING: Counter changed %0d times after pause (may be in-flight instructions)", pause_errors);
      // Don't count as error if it only changed once then stayed stable
      if (pause_errors > 1) begin
        test_errors = test_errors + 1;
      end
    end
    $display("");
    
    // Test 7: Resume Functionality
    $display("━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━");
    $display("TEST 7: Resume Functionality (SW[0] = 1)");
    $display("━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━");
    
    io_sw = 32'h1;  // Set SW[0] = 1 to resume
    $display("  SW[0] = 1 (counter resumed)");
    
    last_counter_value = get_counter_value();
    $display("  Value at resume: 0x%h", last_counter_value);
    
    wait_for_increment(1000, "Resume increment");
    
    current_counter_value = get_counter_value();
    
    if (current_counter_value != last_counter_value) begin
      $display("  ✅ PASS: Counter resumed successfully (0x%h -> 0x%h)",
               last_counter_value, current_counter_value);
    end else begin
      $display("  ❌ FAIL: Counter did not resume");
      test_errors = test_errors + 1;
    end
    
    display_hexleds("After resume");
    $display("");
    
    // Test 8: Memory Address Verification
    $display("━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━");
    $display("TEST 8: Memory-Mapped I/O Addresses");
    $display("━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━");
    
    $display("  Expected memory map (milestone-2):");
    $display("    HEX0-3:  0x1000_2000 - 0x1000_2FFF");
    $display("    HEX4-7:  0x1000_3000 - 0x1000_3FFF");
    $display("    SW:      0x1001_0000 - 0x1001_0FFF");
    $display("");
    
    // For simple counter without SW control, just verify outputs are being written
    // Check that counter continues to change (proves memory writes are working)
    addr_test_errors = 0;
    for (int cycle = 0; cycle < 3; cycle++) begin
      start_value = get_counter_value();
      repeat(500) @(posedge clk);  // Short wait
      end_value = get_counter_value();
      
      $display("  Cycle %0d: Start=0x%h, End=0x%h %s",
               cycle+1, start_value, end_value,
               (end_value != start_value) ? "✓" : "❌");
      
      if (end_value == start_value) begin
        addr_test_errors = addr_test_errors + 1;
      end
    end
    
    if (addr_test_errors == 0) begin
      $display("  ✅ PASS: Memory-mapped I/O working correctly");
    end else begin
      $display("  ❌ FAIL: Memory writes not occurring");
      test_errors = test_errors + 1;
    end
    $display("");
    
    // Test 9: Edge Case Testing
    $display("━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━");
    $display("TEST 9: Edge Cases & Boundary Conditions");
    $display("━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━");
    
    // Check for digit rollovers (e.g., x9 -> y0)
    current_counter_value = get_counter_value();
    ones = decode_7seg(io_hex0);
    tens = decode_7seg(io_hex1);
    
    $display("  Current value: 0x%h (ones=%0d, tens=%0d)", current_counter_value, ones, tens);
    
    // If we're close to a rollover, watch for it
    if (ones == 9) begin
      $display("  Ones digit is 9, watching for rollover to 0...");
      wait_for_increment(5000, "Ones rollover");
      
      new_ones = decode_7seg(io_hex0);
      new_tens = decode_7seg(io_hex1);
      
      if (new_ones == 0 && new_tens == tens + 1) begin
        $display("  ✅ PASS: Ones digit rolled over correctly (9 -> 0, tens incremented)");
      end else if (new_ones == 0 && new_tens == 0 && tens == 9) begin
        $display("  ✅ PASS: Tens digit rolled over correctly (99 -> 00)");
      end else begin
        $display("  ⚠️  Rollover result: ones=%0d, tens=%0d", new_ones, new_tens);
      end
    end else begin
      $display("  ⚠️  Ones digit not at 9, cannot test rollover in this run");
    end
    
    // Verify no glitches in display
    if (all_digits_valid()) begin
      $display("  ✅ PASS: No display glitches detected");
    end else begin
      $display("  ❌ FAIL: Display glitch detected");
      test_errors = test_errors + 1;
    end
    $display("");
    
    // Test 9: Performance Check
    $display("━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━");
    $display("TEST 9: Performance & Timing");
    $display("━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━");
    
    start_cycles = cycle_count;
    start_value = get_counter_value();
    
    // Wait for 3 increments
    for (int i = 0; i < 3; i++) begin
      wait_for_increment(5000, $sformatf("Increment %0d/3", i+1));
    end
    
    elapsed_cycles = cycle_count - start_cycles;
    end_value = get_counter_value();
    
    $display("  Performance metrics:");
    $display("    Cycles elapsed: %0d", elapsed_cycles);
    $display("    Start value: 0x%h", start_value);
    $display("    End value: 0x%h", end_value);
    
    if (end_value != start_value) begin
      $display("  ✅ PASS: Counter incremented (BCD changes detected)");
    end else begin
      $display("  ⚠️  Counter did not change");
    end
    $display("");
    
    // Final summary
    $display("━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━");
    $display("TEST SUMMARY");
    $display("━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━");
    $display("");
    
    display_hexleds("Final State");
    $display("");
    
    if (test_errors == 0) begin
      $display("  ╔══════════════════════════════════════════════════════════════╗");
      $display("  ║  ✅✅✅  ALL TESTS PASSED - HEXLED FULLY FUNCTIONAL  ✅✅✅  ║");
      $display("  ╚══════════════════════════════════════════════════════════════╝");
      $display("");
      $display("  ✓ Display encoding: CORRECT");
      $display("  ✓ Counter logic: WORKING");
      $display("  ✓ Pause/Resume: FUNCTIONAL");
      $display("  ✓ Memory I/O: VERIFIED");
      $display("  ✓ Edge cases: HANDLED");
    end else begin
      $display("  ╔══════════════════════════════════════════════════════════════╗");
      $display("  ║  ❌ %2d TEST(S) FAILED - REVIEW REQUIRED ❌                  ║", test_errors);
      $display("  ╚══════════════════════════════════════════════════════════════╝");
      $display("");
      $display("  Please review the failures above and check:");
      $display("  - counter_v3_fast.hex is loaded correctly");
      $display("  - Memory addresses match milestone-2 spec");
      $display("  - 7-segment encoding table is correct");
    end
    
    $display("");
    $display("  Processor Statistics:");
    $display("    Final PC: 0x%h", pc_commit);
    $display("    Total cycles: %0d", cycle_count);
    $display("    Final counter value: %0d", get_counter_value());
    $display("");
    $display("╔══════════════════════════════════════════════════════════════════╗");
    $display("║                  In-Depth Test Complete                          ║");
    $display("╚══════════════════════════════════════════════════════════════════╝");
    $display("");
    
    $finish;
  end
  
  // Cycle counter
  always @(posedge clk) begin
    if (reset) cycle_count <= cycle_count + 1;
  end

endmodule
